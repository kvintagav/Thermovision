module bufer_line_dual(

);




endmodule

