module xor_value(



)