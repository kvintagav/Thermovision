// megafunction wizard: %Gamma Corrector v11.0%
// GENERATION: DEFERRED
// synthesis translate_off

module gamma (
	clock,
	reset,
	din_ready,
	din_valid,
	din_data,
	din_startofpacket,
	din_endofpacket,
	dout_ready,
	dout_valid,
	dout_data,
	dout_startofpacket,
	dout_endofpacket,
	gamma_lut_0_av_chipselect,
	gamma_lut_0_av_write,
	gamma_lut_0_av_address,
	gamma_lut_0_av_writedata,
	gamma_lut_0_av_readdata,
	gamma_lut_1_av_chipselect,
	gamma_lut_1_av_write,
	gamma_lut_1_av_address,
	gamma_lut_1_av_writedata,
	gamma_lut_1_av_readdata,
	gamma_lut_2_av_chipselect,
	gamma_lut_2_av_write,
	gamma_lut_2_av_address,
	gamma_lut_2_av_writedata,
	gamma_lut_2_av_readdata,
	);
	input		clock;
	input		reset;
	output		din_ready;
	input		din_valid;
	input	[17:0]	din_data;
	input		din_startofpacket;
	input		din_endofpacket;
	input		dout_ready;
	output		dout_valid;
	output	[17:0]	dout_data;
	output		dout_startofpacket;
	output		dout_endofpacket;
	input		gamma_lut_0_av_chipselect;
	input		gamma_lut_0_av_write;
	input	[6:0]	gamma_lut_0_av_address;
	input	[5:0]	gamma_lut_0_av_writedata;
	output	[5:0]	gamma_lut_0_av_readdata;
	input		gamma_lut_1_av_chipselect;
	input		gamma_lut_1_av_write;
	input	[6:0]	gamma_lut_1_av_address;
	input	[5:0]	gamma_lut_1_av_writedata;
	output	[5:0]	gamma_lut_1_av_readdata;
	input		gamma_lut_2_av_chipselect;
	input		gamma_lut_2_av_write;
	input	[6:0]	gamma_lut_2_av_address;
	input	[5:0]	gamma_lut_2_av_writedata;
	output	[5:0]	gamma_lut_2_av_readdata;
endmodule
// synthesis translate_on
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2013 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="alt_vip_gam" version="11.0" >
// Retrieval info: 	<generic name="AUTO_DEVICE_FAMILY" value="Cyclone IV E" />
// Retrieval info: 	<generic name="PARAMETERISATION" value="&lt;gammaParams&gt;&lt;GAM_NAME&gt;MyGammaCorrector&lt;/GAM_NAME&gt;&lt;GAM_CHANNEL_COUNT&gt;3&lt;/GAM_CHANNEL_COUNT&gt;&lt;GAM_CHANNELS_ARE_IN_PAR&gt;true&lt;/GAM_CHANNELS_ARE_IN_PAR&gt;&lt;GAM_BPS&gt;6&lt;/GAM_BPS&gt;&lt;GAM_COMPILE_TIME&gt;false&lt;/GAM_COMPILE_TIME&gt;&lt;GAM_LUT /&gt;&lt;/gammaParams&gt;" />
// Retrieval info: </instance>
