module beaten_pix(

input CLK;
input wire [`ADC_WIDHT-1:0] IN_ADC1;
input wire {`ADC_WIDHT-1:0] IN_ADC2;

output [`ADC_WIDHT-1:0] OUT_ADC1;
output {`ADC_WIDHT-1:0] OUT_ADC2;


);
