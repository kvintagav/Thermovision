// megafunction wizard: %Median Filter 2D v11.0%
// GENERATION: DEFERRED
// synthesis translate_off

module median (
	clock,
	reset,
	din_ready,
	din_valid,
	din_data,
	din_startofpacket,
	din_endofpacket,
	dout_ready,
	dout_valid,
	dout_data,
	dout_startofpacket,
	dout_endofpacket,
	);
	input		clock;
	input		reset;
	output		din_ready;
	input		din_valid;
	input	[13:0]	din_data;
	input		din_startofpacket;
	input		din_endofpacket;
	input		dout_ready;
	output		dout_valid;
	output	[13:0]	dout_data;
	output		dout_startofpacket;
	output		dout_endofpacket;
endmodule
// synthesis translate_on
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2013 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="alt_vip_med" version="11.0" >
// Retrieval info: 	<generic name="AUTO_DEVICE_FAMILY" value="Cyclone IV E" />
// Retrieval info: 	<generic name="PARAMETERISATION" value="&lt;medParams&gt;&lt;MED_NAME&gt;my_mFilter&lt;/MED_NAME&gt;&lt;MED_WIDTH&gt;640&lt;/MED_WIDTH&gt;&lt;MED_HEIGHT&gt;480&lt;/MED_HEIGHT&gt;&lt;MED_FILTER_SIZE&gt;3&lt;/MED_FILTER_SIZE&gt;&lt;MED_BPS&gt;14&lt;/MED_BPS&gt;&lt;MED_CHANNELS_IN_SEQ&gt;1&lt;/MED_CHANNELS_IN_SEQ&gt;&lt;/medParams&gt;" />
// Retrieval info: </instance>
